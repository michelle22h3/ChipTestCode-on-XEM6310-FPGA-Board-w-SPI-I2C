// -------------------------------------------------------------------------------------
// Testbench for FPGA tester top module
// Reference: https://docs.opalkelly.com/display/FPSDK/FrontPanel+HDL+-+Host+Simulation
// -------------------------------------------------------------------------------------

`timescale 1ns/1ps

module FPGATopTestbench();
    
    `include "config.vh"
    `include "func.v"
    
    localparam CLK_PERIOD = 10.0;          // Clock freq = 100MHz
    localparam NO_MASK    = 32'hFFFF_FFFF; // The mask can be set to cover the bits to be change in those 32 bits
    
    //----------------------------------------------------------------
    // Begin okHostInterface simulation user configurable global data
    //----------------------------------------------------------------
    // REQUIRED: # of clocks between blocks of pipe data
    parameter BlockDelayStates = 5;
    // REQUIRED: # of clocks before block transfer before host interface checks for ready (0-255)
    parameter ReadyCheckDelay = 5;
    // REQUIRED: # of clocks after ready is asserted and check that the block transfer begins (0-255)
    parameter PostReadyDelay = 5;
    // REQUIRED: byte (must be even) length of default PipeIn; Integer 0-2^32
    parameter pipeInSize = max(`ACT_IN_BYTES, `WEIGHT_BYTES);  
    // Choose the maximum one
    // REQUIRED: byte (must be even) length of default PipeOut; Integer 0-2^32
    parameter pipeOutSize = `ACT_OUT_BYTES;
    // Size of array for register set commands.
    parameter registerSetSize = 32;
    
    // Pipes
    integer k;
    reg  [7:0]  pipeIn [0:(pipeInSize-1)];
    initial for (k = 0; k<pipeInSize; k = k+1) pipeIn[k] = 8'h00;
    
    reg  [7:0]  pipeOut [0:(pipeOutSize-1)];
    initial for (k = 0; k<pipeOutSize; k = k+1) pipeOut[k] = 8'h00;
    
    // Registers
    reg [31:0] u32Address  [0:(registerSetSize-1)];
    reg [31:0] u32Data     [0:(registerSetSize-1)];
    reg [31:0] u32Count;

    // Golden reference for activation output
    reg [7:0] golden_ref [`ACT_OUT_BYTES-1:0];
    
    
    //----------------------------------------------------------------
    // Host interface connections
    //----------------------------------------------------------------
    wire    [4:0]       okUH;               // Host interface input signals
    wire    [2:0]       okHU;               // Host interface output signals
    wire    [31:0]      okUHU;              // Host interface bidirectional signals
    wire                okAA;               // Host interface bidirectional signal
    reg                 sys_clkp;           // Differential clock signal (positive)
    reg                 sys_clkn;           // Differential clock signal (negative)
    wire    [7:0]       led;                // LED board connections
    // ---------------------------------------------------------------
    // IC chip interface connections
    // ---------------------------------------------------------------
    wire                CLK_100M;           // 100MHz clock generated by FPGA to IC
    wire                rst_n;              // IC chip reset generated by FPGA to IC (active low)
    wire                A_SPI_CLK;          // Activation SPI clock
    wire                A_SPI_MISO;         // Activation SPI RX data
    wire                A_SPI_MOSI;         // Activation SPI TX data
    wire                W_SPI_CLK;          // Weight SPI clock
    wire                W_SPI_MOSI;         // Weight SPI TX data
    wire                Weight_CS_N;        // Weight SPI chip select (active low)
    wire                Activation_CS_N;    // Activation SPI slave chip select (active low)
    wire                chip_start_mapw;    // 2-cycle trigger signal indicating IC start the weight mapping
    wire                chip_start_calc;    // Trigger indicator from FPGA to IC for start calculation
    
    //----------------------------------------------------------------
    // Differential clock signal generation
    //----------------------------------------------------------------
    initial begin
        sys_clkp = 1'b0;
        forever #(CLK_PERIOD / 2)
            sys_clkp = ~sys_clkp;
    end
    always @(*) sys_clkn = ~sys_clkp;
    
    //----------------------------------------------------------------
    // FPGA Top module (Unit Under Test)
    //----------------------------------------------------------------
    FPGATop UUT (
    .okUH               (okUH),             // Host interface input signals
    .okHU               (okHU),             // Host interface output signals
    .okUHU              (okUHU),            // Host interface bidirectional signals
    .okAA               (okAA),             // Host interface bidirectional signal
    .sys_clkn           (sys_clkn),         // System differential clock input (negative)
    .sys_clkp           (sys_clkp),         // System differential clock input (positive)
    .led                (led),              // On board LED pins
    .A_SPI_CLK          (A_SPI_CLK),        // Activation SPI clock
    .A_SPI_MISO         (A_SPI_MISO),       // Output activation RX SPI data (from slave to master)
    .A_SPI_MOSI         (A_SPI_MOSI),       // Input activation TX SPI data (from master to slave)
    .W_SPI_CLK          (W_SPI_CLK),        // Weight SPI clock
    .W_SPI_MOSI         (W_SPI_MOSI),       // Weight TX SPI data (from master to slave)
    .Weight_CS_N        (Weight_CS_N),      // Weight SPI slave chip select (active low)
    .Activation_CS_N    (Activation_CS_N),  // Activation SPI slave chip select (active low)
    .chip_start_mapw    (chip_start_mapw),  // 2-cycle trigger signal indicating IC start the weight mapping
    .chip_start_calc    (chip_start_calc),  // 2-cycle trigger indicating IC start the calculation
    .CLK_100M           (CLK_100M),         // 100MHz clock from FPGA to IC
    .rst_n              (rst_n)             // Chip reset from FPGA to IC (active low)
    );
    
    // ---------------------------------------------------------------
    // Simplified behavior model of chip
    // ---------------------------------------------------------------
    Chip chip (
    .CLK_100M           (CLK_100M),         // 100MHz clock from FPGA to IC
    .rst_n              (rst_n),            // Chip reset from FPGA to IC (active low)
    .chip_start_mapw    (chip_start_mapw),  // 2-cycle trigger signal indicating IC start the weight mapping
    .chip_start_calc    (chip_start_calc),  // 2-cycle indicator to start the calculation
    .A_SPI_CLK          (A_SPI_CLK),        // Activation SPI clock
    .A_SPI_MOSI         (A_SPI_MOSI),       // Activation SPI data from master to slave
    .A_SPI_CS_n         (Activation_CS_N),  // Activation SPI chip select (active low)
    .A_SPI_MISO         (A_SPI_MISO),       // Activation SPI data from slave to master
    .W_SPI_CLK          (W_SPI_CLK),        // Weight SPI clock
    .W_SPI_MOSI         (W_SPI_MOSI),       // Weight SPI data from master to slave
    .W_SPI_CS_n         (Weight_CS_N)       // Weight SPI chip select (active low)
    );
    
    // ---------------------------------------------------------------
    // Handy task to reset the FPGA internal logics
    // ---------------------------------------------------------------
    task reset();
        begin
            // Send software reset
            SetWireInValue(`SW_RST_ADDR, 32'h0000_0001, NO_MASK);
            UpdateWireIns;
            SetWireInValue(`SW_RST_ADDR, 32'h0000_0000, NO_MASK);
            UpdateWireIns;
        end
    endtask
    
    // ---------------------------------------------------------------
    // Handy task to polling over LSB of the specified trigger out
    // ---------------------------------------------------------------
    task polling_trigger_out(input [7:0] trigger_out_addr);
        reg trigger_active;
        begin
            trigger_active = 0;
            while (trigger_active == 0) begin
                UpdateTriggerOuts;
                trigger_active = IsTriggered(trigger_out_addr, 32'h0000_0001);
            end
        end
    endtask
    
    //----------------------------------------------------------------
    // Main testbench (emulate host end behavior)
    //----------------------------------------------------------------
    integer i, error_counts;
    initial begin
        FrontPanelReset;
        reset();
        
        // Read activation input from memory initialization file and send to chip
        $readmemh("act_in.dat", pipeIn);
        WriteToPipeIn(`ACT_IN_DATA_ADDR, `ACT_IN_BYTES);

        // Read weight input from memory initialization file and send to chip
        $readmemh("weight.dat", pipeIn);
        WriteToPipeIn(`WEIGHT_DATA_ADDR, `WEIGHT_BYTES);
        
        // Polling over computation done status
        polling_trigger_out(`CALC_DONE_ADDR);
        $display("[@time = %t]: Host receives computation done from FPGA.", $time);
        
        // Send activation data (maybe dummy) to retrieve the data calculated by chip
        for (i = 0; i < `ACT_IN_BYTES; i = i + 1) begin
            pipeIn[i] = 0; // Send full 0s for dummy data
        end
        WriteToPipeIn(`ACT_IN_DATA_ADDR, `ACT_IN_BYTES);
        
        // Polling over activation output receive status done
        polling_trigger_out(`ACT_OUT_RX_DONE_ADDR);
        $display("[@time = %t]: Host receives activation RX done from FPGA.", $time);
        
        // Read data from activation output pipe and compare against the golden reference
        error_counts = 0;
        $readmemh("golden_ref.dat", golden_ref);
        ReadFromPipeOut(`ACT_OUT_DATA_ADDR, `ACT_OUT_BYTES);
        for (i = 0; i < pipeOutSize; i = i + 1) begin
            $display("[@time = %t]: Host receives calculated outputs from FPGA: %d", $time, pipeOut[i]);
            if (golden_ref[i] != pipeOut[i]) begin
                error_counts = error_counts + 1;
                $display("ERROR: mismatched data golden ref %d vs. calculated %d", golden_ref[i], pipeOut[i]);
            end
        end
        if (error_counts == 0) begin
            $display("Successful. All calculated data matches with the golden reference :-)");
        end
        else begin
            $display("There are %d mismatches", error_counts);
        end

        # 10000
        $finish;
    end
    
    `include "./okSimLib/okHostCalls.v"
    
endmodule
