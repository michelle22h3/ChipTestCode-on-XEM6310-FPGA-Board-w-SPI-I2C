// Address map

// WireIn
`define SW_RST_ADDR 8'h07
`define ITF_SEL_ADDR 8'h08

// WireOut
`define STA_CHIP_ADDR 8'h27

// TriggerIn
`define SPI_CONFIG_ADDR 8'h47

// PipeIn
`define FIFOA_IN_DATA_ADDR 8'h87

`define FIFOB_OUT_DATA_ADDR 8'hA7

// Number of endpoints requiring `okEH`
`define NUM_ENDPOINTS 4




